`include "vunit_defines.svh"
`timescale 1ns/1ns